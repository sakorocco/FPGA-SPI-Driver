`timescale 1ns / 1ps

module SPI_tb(

    );
    
    
endmodule
